module mainProcessor();
endmodule
